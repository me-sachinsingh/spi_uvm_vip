module top;

endmodule